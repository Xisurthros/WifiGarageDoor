PK   ZsUY5/*  rM    cirkitFile.json�ݎ��v�_��������I�����E�@�D�#D#u$�ǎ1���3�JR��UT���t���3�,n�Uk�~Kk����_��l��ճ_��~��LnU2�|,w����o���~����_v����������}�wuYͷ�Y-�"� )�Y�z��b�uV,T5�TR��Y8���0}�p��\�]�Zw�0�߮����yO��Կ4��ŧ�����9�b��~��7�Y��8��y�-t��2�e��h�L¬��81�`�Ȼ&�)1W��^��K�)�b�3-�p��Y����O���Y$����/b���S,>��g���c����O�O����o�L�&2�1W	K}�R/ŧX|���Rq��,)˟�b�)_8�����e,R|�ŧX|�,�����_��q���������s�ɘÒi���e�鸊�*.�A�B�q^˲��EI��크1�[8[8��s�R�5��p�䪗�e/�^b�
��`��� �V�h	аhV��\�R���`!KQ��t�\�R���`9KQ��t�\�R���`QKQ��t�\�R�<�`}�q��V	�l�(�wLo��-�[
��Qy .�H��Ur}L���21D�8��D:������F6\ �.&��`�
�h�L.Q)X�R�H%��`�
�δ\lҰؤa�IQ��t�\lҰؤa�IQ��tpf�>4E���M��`�I��&�M��Q�M���&�M��Q�M���&�M��Q�M��#+FV��E}� (d��.!8.���
��(+Pb�
��`����2��e$�Hb�
��`����2��e$�Hb�
��^���/i��qQGA��2���2O�R'Uϝo�������y{sG����V����5t�ۛ����7F=oo�=ooN=oo>}�FZvºs����_Xy�Y���k�y���~a�9�X��/�?GV�{{�u<+[���+ᇫD��Z�Yj,a�D�L�����_�d���TY�S�\�i�eh�TYP���VQ��W���D��۟�j�,�*[*�t/�:�3M-�*Q�4Q*���no����va��e�4��_��Xg��v��ɝ!&
��MD���=<�qy�:�.�H�u�����Ш��I��d�D�QA�5�I�!d��I�QA�#���[D<*�4�5����L�'�7�xT�i�kQ�G}�%R�����H<*�4�u�����tJq�|ˈG��@��xT����*�
2�v].� �9�	t�*��/�s�4��������I�$d����0�e���u���L$s����x��d���xM@|sR�HZ�Hb���$����)L0s��$ߘf6
n��7&�9V|X�oL9�����S>,�7�������Ih�����[�a�	�GF��	"f%�1���ƴ�Qp{�2�����4��K�)j܄�2
��D�8��c	��j���Xa@|cҚ���%��p{�2���yL_s�%���L_��^���'
>,�7�����c���H�D�HGҸ3i#JG_Ә��[�aI�1}m�s�oL_s|0��$ߘ�6
n��7��9�|X�o��(�=�!ߘ���a�aI�SJ��Ò|c��c}��%����Qp{�? �1}�1��Ò|c��(�=!ߘ���i�aI�1}m�7_���"@�墿��e���p�Ҳ"�o?Di����� QZ���$D�zێK�+!�0�vVb��	���g�M�Q���6���݉�w��I���#���C�(�>N]�?|[����s���q=JW ʫ�t5��޻]9����Lc(5`����r-[ ;��訧ե'�03 =��}2�@8q^��QA�!�3:*ȴ�8q^��QA�!�3:*�tDq⼼���LC�=ftT����ymGG��@{�4� �	ŉ��
2���i�QA�S��Ud�1Ӡ��Lg'�K::*�4�c�AG��)N��stT�i��L��
2]P�8/�� �h���TN0��5��Ò�	�����g����Ie#ie#�e�Z6�\6�^�0��5��Ò|c��(�}fߘl�J�aI�1�l�>3�oL<sM%�$ߘ~6
n���7&���xX�oLE��L���\S	<,�7�����g�����i����S�F��3�`��D5�TK��j����i0|cҚk*��%��ԵQp��4��*���J�a�#+��6
n���7����xX�oL_��L��;�6҉����qg�F:�6���1}�5��Ò|c��(�}fߘ��J�aI�1}m�>3�oL_sM%�$ߘ�6
n���7����xX�oL_��L����\S	<,�7�����g�����k������F��3�`���5�TK��k����ix�0ӐGiQ.�iȣ���iȣ���iȣ��^�4�QZ��!f@�zێK1� �0�vf`�����gC�4�Q���6�x���<
�˫Tg3y�W��fW�t6ӐGy���f�(����LC�e._�毿�ݮ��٪�mr���ϫ]��ݯ�E]�V��vWջ��ݝ��RWQ��@GI�i��<,�A<O�p-tZ���hA�x�a:<��]�E�E&b������9��7D�]��7���f�Jz�R��{�N�J��He���j���u���Te�/�2�Q��2�B�A�5[]��(MM�	3i�zf��E�\Z�>\�j#����N/�̕����E�I�i,�C�����]�i��Yu��ʷ �39��U���(!x1�I�ͬ|�|��M��r��ܛY�='�v��)Ɨ��	������Uw�$荅<#z���l3��W�����vEnBolx���NC����"	�]��%���s���#̔_}��>�u,�Q��n�,p;�w��� O�V��`J�a�yrU�y�\�>�Z�?�*�p}���x�SG3�P(��1V/�c�!⓷���]\<�T1D��:aQ�{���aQ����CX���|�����(���>��!,��^w�S��CXC���s�NӮ�_qL�$8_���!��!z,̹xȣ��{��:aQ�cO��CX���|ɉ���(����!,��-�[<��BR��0	I��$8��؍7�G2�9'η��xǅ�iBe�E�1�
�,�l�P�`�>q)����A�DB�"DKB
Є\sl0 �% �(}��R.e�5�2\���g�-�Ї\Sk0 �% �(}��R.Y�5�2\&�62A+E0�3��	Z,r]���r����(�DH-  �6�`@�Z@CrQ6��P�A����L�:��5-�P�`�>Gm)��\�I�.�(}��`@�| �N�`@� �(}N�R.��u�2\"���r-�88��g���C�H���uo2\"���N-��\gf0 �% �(}��R.��u]2\Ǉ`�>Wi)��*�:*�.Sw��	�p@��a�\/e0 �4 �(}^�R.U��I2\����-�P�\d0 �%�
�(}��;K�w���%�;��.Β���� �f����1��Yr��qh�V�{ve��(����CܗE�u�L�,����j�����Z`�|�� ��k��._{�<�}Y�����?\g�t:[/����tYr����l���N%�)��Z/?�YU���&��~����:���د�ټ�cf��>�
-�v+l��ͱ�m�lSe�*�X���6W���7({��whk�9�R�ɘ ]*�9����7t!����N����g��mn���;��}x��F�n��*C�o�F��PK�0�ugGA>���%	����;��;﫸ܺS� 9�z�y,>��`]���ݱx�����T�Q�x)q/��K�{);_��K�|I����Ƚ��/���|)t/��%e��z={Qʫ�r;[��KWZf*\Ƌ���8�Y����X'�Ϊ����h�g�=��h�����BL>�i�֛���L'����Rkv�g<�����Ci��q�ջ����V�q���~c��Ehzpح6��mS~�?۫�ɯ�����sm������:1��~�q�&��vY������w?�����~�ݮ�χծ�&�����S�yX����Κ1���f�i�CU.w��7�o�{O��2i��huXmM�ܩ4��m���c�i��DY�&��3]l��D�D�E�<��4+�"N��,����"]�q���g���r�8��iq:�l�͡<%69��b�[��3�wZ��}*�i����yrsz�G;��ά+[�S U�5�l����� ?_N.F����~@Z��}-͒�S���,Ӥ�Aq�8�=�{��s3�T��|��)�<�FOѲ�j��8G�IK��ܕ��Az"#��#%�4{��j���5�(2Oo��ڙr�p|,�cu���P��?׻��Q7��n=���S��F�qX(������SG<?�w�r��T��z��Am�Z�^���|�,���w��5���ꗏ���Gi'�y�vSG7fߧ�0~lv�MU�'�%�\�.���*�� ��D�yr�b�$ab���n�E��y��XZ���3���_���ԯ/��j�`�����E���C���4�?�ݘ(�М�w�����_�:�vx(
�ę)�B�E�߶�z���$\m?o��yn�<�%�|�[���M��>�*�Q�?�?����N?��s�g�sfٿ<|�׻o~\~�m���W�k�}��E��ԌY�>�9���Ȏ�Q����4��e�q�IR&A��eg�|��͇���|��j��)m��SBw�p�{aPm�YM�˿��.��T��%շ�mY8�:*o����#F�M�<���P?v�����*�T�C��V��[�/��2�sU-R}T�.j����ie畋q�x,υ|؄�o��o�:���}0;	�:�ݘ����NudG�H��\CF]��|a��yl��i�ٵsa�6�n��ӨX4ˣ���,���xYQ�(ҩY+ބc�q�s�EffLr�ʹ.��j��������>�H⣾|,_3��>gb�͛����&5˖�,&m�|����K�B6MmwԿ]���˰VG/��ۧ��]}8�������ձ���'��������Ofh��'��������j�}u�$�l��M�	�W>>�ڕ�z5�`�0��{|�5~���\������<|<���������|g/�t|d����w��:�/�m��`>�gL��"�ne�����Vv��Շ/�'_Lu5J%������W��R&ba����kk�0��,��O���ZQ�i�X�����w����sm��5�K'�KǓ��t��vɵ����)���jp�y���O��x3���Wf,&y�v�^) ��� �:�.��[����]�� 7*�Ow2�U�x[�Ev���k}��Q"sy��a��m��y�'���'q�$.���������m�w�b�Y>V�8�X�V|��I�g!žW�oL/]��5jt;��25z�
��ɶ��������I��V�Ө��4�������H,O���Q��E���Z�ƒ��R�X%p�^����<ԻU���2��?��������<��o���?ԟ�Ї/�/�PK
   ZsUY5/*  rM                  cirkitFile.jsonPK      =   E    